-- Test file for "God-Tier" static analysis rules
-- This file intentionally contains violations to test the advanced rules

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- =============================================================================
-- Test 1: Hardware Trojan Detection (Security Analysis)
-- =============================================================================

entity trojan_test is
    port (
        clk        : in  std_logic;
        rst_n      : in  std_logic;
        counter    : in  std_logic_vector(31 downto 0);
        data_in    : in  std_logic_vector(31 downto 0);
        secret_out : out std_logic;
        normal_out : out std_logic_vector(7 downto 0)
    );
end entity trojan_test;

architecture rtl of trojan_test is
    signal trigger : std_logic;
begin
    -- TROJAN PATTERN: Magic number comparison driving output
    -- This should trigger multiple security rules:
    -- 1. magic_number_comparison (DEADBEEF is a known magic number)
    -- 2. trigger_drives_output (comparison drives output port)
    trojan_proc: process(clk, rst_n)
    begin
        if rst_n = '0' then
            secret_out <= '0';
        elsif rising_edge(clk) then
            -- This is a classic trojan trigger pattern!
            if counter = X"DEADBEEF" then
                secret_out <= '1';  -- Kill switch activates
            end if;
        end if;
    end process;

    -- Another suspicious pattern: large literal comparison
    -- Should trigger large_literal_comparison
    counter_check: process(clk)
    begin
        if rising_edge(clk) then
            if counter = X"CAFEBABE" then
                trigger <= '1';
            end if;
        end if;
    end process;
end architecture rtl;

-- =============================================================================
-- Test 2: Reset Domain Crossing (RDC Analysis)
-- =============================================================================

entity rdc_test is
    port (
        clk_a    : in  std_logic;
        clk_b    : in  std_logic;
        rst_async: in  std_logic;
        data_a   : in  std_logic_vector(7 downto 0);
        data_b   : out std_logic_vector(7 downto 0)
    );
end entity rdc_test;

architecture rtl of rdc_test is
    signal reg_a : std_logic_vector(7 downto 0);
    signal reg_b : std_logic_vector(7 downto 0);
    -- Combinationally generated reset (BAD!)
    signal gen_rst : std_logic;
begin
    -- BAD: Same reset used in two different clock domains
    -- Should trigger reset_crosses_domains
    domain_a: process(clk_a, rst_async)
    begin
        if rst_async = '1' then
            reg_a <= (others => '0');
        elsif rising_edge(clk_a) then
            reg_a <= data_a;
        end if;
    end process;

    domain_b: process(clk_b, rst_async)
    begin
        if rst_async = '1' then
            reg_b <= (others => '0');
        elsif rising_edge(clk_b) then
            reg_b <= reg_a;
            data_b <= reg_b;
        end if;
    end process;

    -- BAD: Reset generated by combinational logic
    -- Should trigger combinational_reset_gen
    gen_rst <= rst_async and data_a(0);
end architecture rtl;

-- =============================================================================
-- Test 3: Combinational Loop Detection
-- =============================================================================

entity loop_test is
    port (
        a_in  : in  std_logic;
        b_in  : in  std_logic;
        c_out : out std_logic
    );
end entity loop_test;

architecture rtl of loop_test is
    signal x, y, z : std_logic;
begin
    -- Direct combinational loop: x depends on itself
    -- Should trigger direct_combinational_loop
    x <= x and a_in;

    -- Two-stage loop: y -> z -> y
    -- Should trigger two_stage_loop
    y <= z and a_in;
    z <= y or b_in;

    c_out <= x xor y;
end architecture rtl;

-- =============================================================================
-- Test 4: Power Vampire (Operand Isolation)
-- =============================================================================

entity power_test is
    port (
        clk      : in  std_logic;
        rst      : in  std_logic;
        enable   : in  std_logic;
        a        : in  unsigned(15 downto 0);
        b        : in  unsigned(15 downto 0);
        result   : out unsigned(31 downto 0);
        quotient : out unsigned(15 downto 0)
    );
end entity power_test;

architecture rtl of power_test is
    signal mult_result : unsigned(31 downto 0);
    signal div_result  : unsigned(15 downto 0);
begin
    -- POWER VAMPIRE: Unguarded multiplication
    -- Should trigger unguarded_multiplication
    -- This multiplier runs EVERY clock cycle even when result isn't used!
    mult_proc: process(clk)
    begin
        if rising_edge(clk) then
            mult_result <= a * b;  -- BAD: No enable guard
            result <= mult_result;
        end if;
    end process;

    -- WORSE: Unguarded division
    -- Should trigger unguarded_division (ERROR severity)
    div_proc: process(clk)
    begin
        if rising_edge(clk) then
            div_result <= a / b;  -- VERY BAD: Division runs every cycle!
            quotient <= div_result;
        end if;
    end process;

    -- GOOD PATTERN (for comparison): Guarded multiplication
    -- This should NOT trigger violations
    good_proc: process(clk)
    begin
        if rising_edge(clk) then
            if enable = '1' then
                -- Multiplier only active when enabled
                result <= a * b;
            end if;
        end if;
    end process;
end architecture rtl;

-- =============================================================================
-- Test 5: Combined Issues (Multiple God-Tier Rules)
-- =============================================================================

entity combined_test is
    port (
        clk     : in  std_logic;
        rst     : in  std_logic;
        trigger : in  std_logic_vector(63 downto 0);
        payload : out std_logic
    );
end entity combined_test;

architecture rtl of combined_test is
    signal internal : std_logic;
    signal counter  : unsigned(31 downto 0);
begin
    -- Multiple suspicious comparisons in same process
    -- Should trigger multi_trigger_process
    suspicious_proc: process(clk, rst)
    begin
        if rst = '1' then
            internal <= '0';
            payload <= '0';
        elsif rising_edge(clk) then
            -- Multiple magic number checks = very suspicious!
            if trigger = X"DEADC0DE12345678" then
                internal <= '1';
            end if;
            if counter = X"BAADF00D" then
                internal <= '1';
            end if;
            if trigger(31 downto 0) = X"FEEDFACE" then
                payload <= internal;
            end if;
        end if;
    end process;
end architecture rtl;
