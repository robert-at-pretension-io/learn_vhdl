library ieee;
use ieee.std_logic_1164.all;

entity demo_tb is
  port (
    clk : in std_logic
  );
end demo_tb;

architecture rtl of demo_tb is
begin
  null;
end rtl;

entity dut is
  port (
    a : in std_logic
  );
end dut;

architecture tb of dut is
begin
  null;
end tb;
