-- Your test VHDL code goes here
-- Start simple and build up!

-- Example: uncomment when you add entity support
-- entity counter is
-- end entity counter;
