package test is
    type state_type is (IDLE, RUN, DONE);
end package test;
