function foo return integer is
begin
    shift_reg(i) <= shift_reg(i);
end;
