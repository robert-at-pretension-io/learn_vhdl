configuration cfg_missing of missing_entity is
end configuration cfg_missing;
