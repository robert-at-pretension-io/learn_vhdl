function foo return integer is
begin
end;
