function foo return integer is
begin
    uniform(seed1, seed2, result);
end;
