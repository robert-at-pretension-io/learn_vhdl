-- minimal function body
function foo return integer is
begin
end function;
