function foo return integer is
begin
    bar(x);
end;
