function foo return integer is
begin
    for i in 0 to 10 loop
        x := x + 1;
    end loop;
end;
