function foo return integer is
begin
    bar(123);
end;
