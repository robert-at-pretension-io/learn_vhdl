function foo return integer is
begin
    bar;
end;
