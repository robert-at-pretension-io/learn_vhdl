function foo return integer is
begin
    shift_reg(i+1) <= shift_reg(i);
end;
