function foo return integer is
begin
    while x > 1 loop
        x := x + 1;
    end loop;
end;
