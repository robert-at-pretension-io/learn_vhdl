package phys_pkg is
  type time_t is range 0 to 1 units
    ns;
    us = 1000 ns;
  end units;
end package;
