function foo return integer;
