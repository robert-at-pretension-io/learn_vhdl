package body test is
    function foo return integer is
    begin
        return 1;
    end function foo;
end package body test;
