package subprograms_rules is
  function bad_fn(a : out integer) return integer;
  procedure bad_proc(b : buffer integer);
end subprograms_rules;
