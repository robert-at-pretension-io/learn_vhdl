-- Minimal test for debugging
package test is
    function log2(n : positive) return natural;
end package test;
