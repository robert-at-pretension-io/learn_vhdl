function foo return integer is
begin
    while i < 8 loop
        x := 1;
    end loop;
end;
